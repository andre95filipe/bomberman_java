10.227.156.4
6666